library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use work.new_types.all;

entity spectra_memory is

end spectra_memory;

architecture Behavioral of spectra_memory is

begin


end Behavioral;
